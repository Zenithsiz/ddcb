pBAV       �� ��# Z  d@  ����	x��@�  ��������x��@�  ��������d��-�  ��������F��@�  ��������_��-�  ��������i��F�  ��������f��@�  ��������2��F�  ��������  �� �  ��������	s��@�  ��������\��@�  ��������N��F�  ��������\��@�  ��������N��(�  ��������n��@�  ��������`��@�  ��������  �� �  ����������@�  ��������U��-�  ��������n��@�  ��������n��@�  ��������d��K�  ��������i��@�  ��������F��@�  ��������  �� �  ��������n��@�  ��������s��@�  ��������P��@�  ��������\��@�  ��������Z��@�  ��������_��@�  ��������F��@�  ��������A��F�  ��������N��-�  ��������  �� �  ��������Z��@�  ��������d��-�  ��������A��@�  ��������Z��@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  n@/ ##      ��� ��   � � � �  n@2 &&      ��� ��   � � � �  PP, **      �����_   � � � �  UP;{..      ��ʀCN   � � � �  x@D 11      ��� ��   � � � �  n> --      ��� ��   � � � �  n(> ))      ��� ��   � � � �  X-Hr;;      ��� k�   � � � �   A@& &&      ��� ��   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   n@8o x    ��݀�O  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@=t x      �����O 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@U~ x      �����_ 
 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@Yz x      ��܀GP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@=v x    �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@Nt x    ��܀GQ  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@Nj x    ��܀GQ  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n@- $$      ��� ��	  � � � �  dP!       �����_	  � � � �  @E 44      ��� ��	  � � � �  i2b JJ      ��� ��	  � � � �  i(n MM      ��� ��	  � � � �  xF^??      ��� ��	  � � � �  Z-        ��� ��	  � � � �  n@R ::      ��� ��	  � � � �  d@J 44      ��� ��	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �  n.| $      ��܀JQ
  � � � �  n@.|%)      ��܀JQ
  � � � �  nF.|*x      ��܀JQ
  � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �               �����_
   � � � �  nF~ =      ��݀EP  � � � �  n@F~>D      ��݀EP  � � � �  nFF~Ex      ��݀EP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  d@Nj x    ���GP  � � � �  n@Zt x    ���GP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@Z` x    ���GP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n@:t x      ����GP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@^t x      ����JP  � � � �  Z@Rj x      ����GP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   x@/ ##      ��� ��  � � � �  PP, **      �����_  � � � �  UP;{..      ��ʀCN  � � � �  x@D 11      ��� ��  � � � �  xF: --      ��� ��  � � � �  xP: ))      ��� ��  � � � �  X-Hr;;      ��� k�  � � � �  U@( &&      ��� ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@=t x      �����O 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n@:t x    ����EP  � � � �   <@8o x    �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@^t x      ��̀R  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@=v x    ��܀�O  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n@a{ x      ��ʀ�M  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@aq x      ��ʀ�M  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  x@E  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   x@/ ##      ��� ��  � � � �  n@0 &&      ��� ��  � � � �  KP( **      �����_  � � � �  FP7{..      ��ʀM  � � � �  x@@ 11      ��� >�  � � � �  n> --      ��� ��  � � � �  n(> ))      ��� ��  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  njw]]      �����_  � � � �  <ec]]      �����_  � � � �  n(kw^^      �����_  � � � �  <(fc^^      �����_  � � � �  n2lw__      �����_  � � � �  <2gc__      �����_  � � � �  n@mw``      �����_  � � � �  <@hc``      �����_  � � � �  nFnwaa      �����_  � � � �  <Ficaa      �����_  � � � �  nPowbb      �����_  � � � �  <Pjcbb      �����_  � � � �  nZpwcc      �����_  � � � �  <Zkccc      �����_  � � � �  ndqwdd      �����_  � � � �  <dlcdd      �����_  � � � �   d@:q x      �����O  � � � �   d@Do x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@Rz x     ��̑
P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@b{ x      ��ݪEP  � � � �  d2nq x      ��ݪEP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   n@d} x    �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  n@P  x      �����_   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  n@U{ x      ��ʥ�P!  � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �               �����_!   � � � �  n@U~ x    �����O# 
 � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �               �����_#   � � � �  n@U{ x      ��ʑ
M$  � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �               �����_$   � � � �  n@Yv x      ����M%  � � � �  <@Ab x      ����M%  � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �               �����_%   � � � �   nFU{99      �����_&  � � � �   n2U{EE      �����_&  � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �               �����_&   � � � �   � 
r � jL�X�rZ�b � n � JXP�� D �N r` ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                