pBAV       �x ��   Z@  ������@�  ��������n��@�  ����������@�  ����������@�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  �������� @=} x      ������   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  o@A  M      �����  � � � �  x@T NV      �����  � � � �  d@T Wl      �����  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @< $$      �����  � � � �   n@& &&      �����_  � � � �  P@& &&      �����_  � � � �   @+z**      ����%�  � � � �   @/z..      ����e�  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  H  x      �����_  � � � �  ~H
 x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @?} x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   
�
f	� ���T                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              