pBAV       P ��   d@  ����U��@�  ��������z��@�  ��������z��@�  ��������i��@�  ��������v��@�  ��������i��@�  ��������K��@�  ��������z��@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  6`  x      �����_   � � � �   Jl2 x      �����_   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  @9  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  r  x      �����_  � � � �   ~r2 x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   Z(<        �����_  � � � �  d<2       �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   T 0S      �����_  � � � �   ~S 0S      �����_  � � � �   d6x Tx      �����_  � � � �  P6x Tx      �����_  � � � �   6  /      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  x $x      �����_  � � � �  ^ ##      �����_  � � � �   P@ "      �����_  � � � �  F@ "      �����_  � � � �  "       �����_  � � � �          �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   d@H  x      �����_  � � � �  Z@H  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @T  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   ��
�� ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              