pBAV       � �� � ] n@  ������@�  ����������@�  ����������@�  ����������@�  ����������@�  ����������@�  ����������@�  ����������@�  ��������s��@�  ��������s��@�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  �������� @` <<      �����_   � � � �  @e ==      �����_   � � � �  @P >>      �����_   � � � �  @c ??      �����_  	 � � � �  @d @@      �����_   � � � �  d@_ AA      �����_  
 � � � �  d@h BB      �����_  
 � � � �  U@e CC      �����_   � � � �  T@h DD      �����_   � � � �  @h EE      �����_   � � � �  @v FF      �����_   � � � �  d@r GG      �����_   � � � �  @p HH      �����_   � � � �  i@y II      �����_  # � � � �  @n JJ      �����_  $ � � � �    @` KK      �����_   � � � �  s@` <<      �����_  � � � �  l@a ==      �����_  � � � �  x@b >>      �����_  � � � �  p@c ??      �����_  � � � �  p@d @@      �����_  � � � �  i@c AA      �����_  � � � �  x@f BB      �����_  � � � �  z@g CC      �����_  � � � �  n@h DD      �����_  � � � �  u@i EE      �����_  � � � �  @v FF      �����_  � � � �  u@n GG      �����_  � � � �  p@l HH      �����_  � � � �  n@m II      �����_  � � � �  i@n JJ      �����_  � � � �  w@o KK      �����_  � � � �  v@` <<      �����_  � � � �  @d ==      �����_  � � � �  s@b >>      �����_  � � � �  s@f ??      �����_  � � � �  x@n @@      �����_  � � � �  o@e AA      �����_  � � � �  o@f BB      �����_   � � � �  o@g CC      �����_ ! � � � �  @h DD      �����_ " � � � �    @h EE      �����_ " � � � �    @h FF      �����_ " � � � �    @h GG      �����_ " � � � �    @h HH      �����_ " � � � �    @h II      �����_ " � � � �    @h JJ      �����_ " � � � �    @h KK      �����_ " � � � �  n@` <<      �����_ % � � � �    @d ==      �����_ % � � � �    @b >>      �����_ % � � � �    @i ??      �����_ % � � � �    @n @@      �����_ % � � � �    @e AA      �����_ % � � � �    @f BB      �����_ % � � � �    @g CC      �����_ % � � � �    @h DD      �����_ % � � � �    @h EE      �����_ % � � � �    @h FF      �����_ % � � � �    @h GG      �����_ % � � � �    @h HH      �����_ % � � � �    @h II      �����_ % � � � �    @h JJ      �����_ % � � � �    @h KK      �����_ % � � � �   @l <<      �����_  � � � �   @a ==      �����_  � � � �  z@n >>      �����_ & � � � �  @c ??      �����_ ' � � � �   `@d @@      �����_ ( � � � �    @i AA      �����_  � � � �  l@_ BB      �����_ ) � � � �    @s CC      �����_  � � � �  x@t DD      �����_ * � � � �    @t EE      �����_  � � � �    @t FF      �����_  � � � �    @t GG      �����_  � � � �    @t HH      �����_  � � � �    @t II      �����_  � � � �    @t JJ      �����_  � � � �    @t KK      �����_  � � � �    @` <<      �����_  � � � �    @a ==      �����_  � � � �  @b >>      �����_ + � � � �  l@c ??      �����_ , � � � �  u@d @@      �����_ - � � � �  d@e AA      �����_ . � � � �  \@Z BB      �����_ / � � � �    @f CC      �����_  � � � �  @g DD      �����_ 0 � � � �  u@f EE      �����_ 1 � � � �  b@j FF      �����_ 2 � � � �  x@d GG      �����_ 3 � � � �  z@p HH      �����_ 4 � � � �    @z II      �����_  � � � �  @n JJ      �����_ 5 � � � �  @s KK      �����_ 6 � � � �  s@` <<      �����_ 7 � � � �  @a ==      �����_ 8 � � � �  h@b >>      �����_ 9 � � � �  s@c ??      �����_ : � � � �  }@p @@      �����_ ; � � � �  {@e AA      �����_ < � � � �  x@P BB      �����_ = � � � �  x@] CC      �����_ = � � � �    @V DD      �����_  � � � �  p@] EE      �����_ > � � � �  }@n FF      �����_ > � � � �  z@s GG      �����_ ? � � � �  z@l HH      �����_ @ � � � �    @w II      �����_  � � � �  @z JJ      �����_ A � � � �  @{ KK      �����_ B � � � �  r@\ <<      �����_ C � � � �    @c ==      �����_  � � � �    @b >>      �����_  � � � �    @c ??      �����_  � � � �  @i @@      �����_ D � � � �    @^ AA      �����_  � � � �    @f BB      �����_  � � � �  K@T CC      �����_ E � � � �  r@d DD      �����_ F � � � �    @j EE      �����_  � � � �    @i FF      �����_  � � � �    @_ GG      �����_  � � � �    @k HH      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �    @T <<      �����_  � � � �  @U ==      �����_ G � � � �  d@V >>      �����_ H � � � �  v@W ??      �����_ I � � � �  }@X @@      �����_ J � � � �  }@Y AA      �����_ K � � � �    @Z BB      �����_  � � � �    @g CC      �����_  � � � �  t@[ DD      �����_ L � � � �    @g EE      �����_  � � � �    @] FF      �����_  � � � �  d@W*GG      �����_ M � � � �  @_ HH      �����_ N � � � �  n@_ II      �����_ O � � � �  }@n JJ      �����_ P � � � �    @o KK      �����_  � � � �  @` <<      �����_	 Q � � � �    @U ==      �����_	  � � � �  k@> >>      �����_	 R � � � �    @W ??      �����_	  � � � �    @X @@      �����_	  � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �               �����_	   � � � �   P@T <<      �����_
 U � � � �   d@U ==      �����_
 T � � � �   x@b >>      �����_
 S � � � �   n@U ??      �����_
 V � � � �   n@] @@      �����_
 V � � � �  U@Y AA      �����_
 W � � � �  _@W BB      �����_
 X � � � �  _@P CC      �����_
 Y � � � �  Z@L DD      �����_
 Z � � � �  Z@T EE      �����_
 Z � � � �   d@b FF      �����_
 [ � � � �  d@X GG      �����_
 \ � � � �  n@W HH      �����_
 ] � � � �   @n II      �����O
 ] � � � �   n@} JJ      �����_
  � � � �               �����_
   � � � �   � � D $ � X � N N������ �f� lT (HN��� Z 
�� PD>V PD <�� Zb��� v ��:�R�� �l��> �0� � N �� � X� � ��>
& 0 � � .h t ` �|                                                                                                                                                                                                                                                                                                                                    