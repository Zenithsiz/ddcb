pBAV        O ��  	 Z@  ����t��@�  ��������|��@�  ��������x��@�  ����������@�  ��������|��@�  ��������|��@�  ��������x��@�  ��������x��@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  �������� @L  x    ����IV   � � � �  @X
 x    ����IV   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �  @@  <    �����R  � � � �  @J =x    ��˞�U  � � � �  @4 <    �����R  � � � �  @>=x    ��˞�U  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @C  x    ��܀�O  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @-  x      ����P  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   @Q  x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @9  x      ��ݙN\  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @Q  x      ��ɒHP  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �  @H  x      ����N 	 � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   
P����($\                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            