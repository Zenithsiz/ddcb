pBAV        p ��   n@  ������@�  ����������@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  P@T <<      �����_   � � � �   d@U ==      �����_   � � � �   x@b >>      �����_   � � � �   n@U ??      �����_   � � � �   n@] @@      �����_   � � � �  _@T AA      �����_   � � � �  _@Z BB      �����_   � � � �   x@Y CC      �����_   � � � �  i@Z DD      �����_   � � � �  n@T EE      �����_   � � � �  @U FF      �����_   � � � �  @f GG      �����_   � � � �  n@R HH      �����_  
 � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   U@L <<      �����_  � � � �   i@I ==      �����_  � � � �  d@L >>      �����_  � � � �  x@L ??      �����_  � � � �  x@N @@      �����_  � � � �  @X AA      �����_  � � � �  d@N BB      �����_  � � � �  @b CC      �����_  � � � �  x@F DD      �����_  � � � �  x@U EE      �����_  � � � �  n@J FF      �����_  � � � �  j@S GG      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   � 0 & � � ��J`<�	�	* 
xz�
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  