pBAV       �� �� &  Z@  ����d��@�  ��������u��@�  ��������s��@�  ��������d��@�  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  �� �  ��������  @$ $$      �����_   � � � �   @* **      �����_   � � � �   @. ..      �����_   � � � �   n@& &&      �����_   � � � �   @C ,,      �����_   � � � �  @$ 00      �����_   � � � �  @* 66      �����_   � � � �  @. ::      �����_   � � � �  @& 22      �����_   � � � �  @$       �����_   � � � �  @*       �����_   � � � �  @. ""      �����_   � � � �  @&       �����_   � � � �               �����_    � � � �               �����_    � � � �               �����_    � � � �   TAn ;    �����_  � � � �   xT5n )    �����_  � � � �   T5n*;    ����(N  � � � �   dTen<x      �����_  � � � �  dTed<x      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   TWP==      �����_  � � � �   V
>>      �����_  � � � �   d@V >>      �����_  � � � �   n~V
>>      �����_  � � � �   @K ??      �����_ 	 � � � �   @Y AA      �����_ 
 � � � �   @X @@      �����_  � � � �   @Z BB      �����_  � � � �   @[ CC      �����_  � � � �   @\ DD      �����_  � � � �   @] EE      �����_  � � � �   @^ FF      �����_  � � � �   @_ GG      �����_  � � � �   @` HH      �����_  � � � �   @a II      �����_  � � � �   @b JJ      �����_  � � � �   Tl;;      �����_  � � � �    T^;;      �����_  � � � �    Sl::      �����_  � � � �   S^::      �����_  � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �               �����_   � � � �   � �x���J�� PFL`<���>�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    